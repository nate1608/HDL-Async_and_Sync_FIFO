`timescale 1ns / 1ps

module control(
    input clk,
    input [3:0] wr_ptr, rd_ptr,
    output reg wr_en, rd_en
    );
    
endmodule
